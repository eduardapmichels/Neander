library verilog;
use verilog.vl_types.all;
entity runstep_vlg_vec_tst is
end runstep_vlg_vec_tst;
