library verilog;
use verilog.vl_types.all;
entity CONT3b_vlg_vec_tst is
end CONT3b_vlg_vec_tst;
