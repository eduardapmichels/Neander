library verilog;
use verilog.vl_types.all;
entity DECOD_vlg_vec_tst is
end DECOD_vlg_vec_tst;
