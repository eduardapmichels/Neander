library verilog;
use verilog.vl_types.all;
entity UnidadeControle_vlg_vec_tst is
end UnidadeControle_vlg_vec_tst;
