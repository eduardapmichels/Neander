library verilog;
use verilog.vl_types.all;
entity DECOD3b8b_vlg_vec_tst is
end DECOD3b8b_vlg_vec_tst;
