library verilog;
use verilog.vl_types.all;
entity RUNSTEPmode_vlg_check_tst is
    port(
        clkclk          : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end RUNSTEPmode_vlg_check_tst;
