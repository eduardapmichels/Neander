library verilog;
use verilog.vl_types.all;
entity LAB09_vlg_vec_tst is
end LAB09_vlg_vec_tst;
