library verilog;
use verilog.vl_types.all;
entity DECOD4b16b_vlg_vec_tst is
end DECOD4b16b_vlg_vec_tst;
