library verilog;
use verilog.vl_types.all;
entity teste_dec_cod_vlg_vec_tst is
end teste_dec_cod_vlg_vec_tst;
