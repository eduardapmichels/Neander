library verilog;
use verilog.vl_types.all;
entity CODULA8b3b_vlg_vec_tst is
end CODULA8b3b_vlg_vec_tst;
