library verilog;
use verilog.vl_types.all;
entity TEMPORIZADOR_vlg_vec_tst is
end TEMPORIZADOR_vlg_vec_tst;
