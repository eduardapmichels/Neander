library verilog;
use verilog.vl_types.all;
entity RUNSTEPmode_vlg_vec_tst is
end RUNSTEPmode_vlg_vec_tst;
