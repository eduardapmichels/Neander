library verilog;
use verilog.vl_types.all;
entity register8b_vlg_vec_tst is
end register8b_vlg_vec_tst;
