library verilog;
use verilog.vl_types.all;
entity SpecReg8b_vlg_vec_tst is
end SpecReg8b_vlg_vec_tst;
